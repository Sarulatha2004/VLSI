module buffer(input in,input ctrl, output out);
buf(out,in);
endmodule
