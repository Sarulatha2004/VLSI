module not_gate(a,o);
input a;
output o;
assign o=~a;
endmodule
