module buffer(input in,input ctrl, output out);
bufif1(out,in,ctrl);
endmodule
