module nand_gate(a,b,o);
input a,b;
output o;
nand g1(o,a,b);
endmodule
