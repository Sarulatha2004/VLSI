module and_gate(a,b,o);
input a,b;
output o;
and g1(o,a,b);
endmodule
