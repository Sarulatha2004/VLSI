module buffer(input in,input ctrl, output out);
bufif0(out,in,ctrl);
endmodule
