module tb_dff_blocking;                                                                                                                                       reg d, clk;                                                                                                                                                 wire q;                                                                                                                                                                                                                                                                                                                 dff_blocking uut(d, clk, q);                                                                                                                                                                                                                                                                                            initial begin                                                                                                                                                 $monitor($time, " clk=%b d=%b q=%b", clk, d, q);
    clk = 0; d = 0;                                                                                                                                             #5 d = 1;                                                                                                                                                   #10 d = 0;
    #20 $finish;                                                                                                                                              end                                                                                                                                                                                                                                                                                                                     always #5 clk = ~clk;                                                                                                                                     endmodule  
