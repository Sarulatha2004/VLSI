module tb_2bit_comp;
reg [1:0]a,b;
wire eq,lt,gt;
comp_2bit uut( .a(a), .b(b), .eq(eq), .lt(lt), .gt(gt));
initial begin
	$dumpfile("2bit_comp_wave.vcd");
	$dumpvars(0, tb_2bit_comp);
	$display("            2 bit comparator               ");
	$display("-------------------------------------------");
	$display("  A       B     |    A>B   A==B    A<B");
	$monitor(" %b %b     %b %b    |     %b     %b       %b",a[1],a[0],b[1],b[0],gt,eq,lt);
        a[1]=0; a[0]=0; b[1]=0; b[0]=0; #10;
        a[1]=0; a[0]=0; b[1]=0; b[0]=1; #10;
        a[1]=0; a[0]=0; b[1]=1; b[0]=0; #10;
        a[1]=0; a[0]=0; b[1]=1; b[0]=1; #10;
        a[1]=0; a[0]=1; b[1]=0; b[0]=0; #10;
        a[1]=0; a[0]=1; b[1]=0; b[0]=1; #10;
        a[1]=0; a[0]=1; b[1]=1; b[0]=0; #10;
        a[1]=0; a[0]=1; b[1]=1; b[0]=1; #10;
        a[1]=1; a[0]=0; b[1]=0; b[0]=0; #10;
        a[1]=1; a[0]=0; b[1]=0; b[0]=1; #10;
        a[1]=1; a[0]=0; b[1]=1; b[0]=0; #10;
        a[1]=1; a[0]=0; b[1]=1; b[0]=1; #10;
        a[1]=1; a[0]=1; b[1]=0; b[0]=0; #10;
        a[1]=1; a[0]=1; b[1]=0; b[0]=1; #10;
        a[1]=1; a[0]=1; b[1]=1; b[0]=0; #10;
        a[1]=1; a[0]=1; b[1]=1; b[0]=1; #10;

$finish;
end
endmodule
