module or_gate(a,b,o);
input a,b;
output o;
or g1(o,a,b);
endmodule

